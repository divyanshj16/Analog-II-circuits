*Differentiator Using OP_AMP
X1 0 3 5 6 4 ua741
R1 1 2 1k
C1 2 3 10n
R2 3 4 10k
C2 3 4 100pf
Vcc 5 0 dc 12v
Vee 0 6 dc 12v
Vin 1 0 pulse(0v 2v 0ms 0ms 0ms 0.1ms .2ms)
.include ua741
.tran .4us 6ms 4ms .001ms
.probe
.end

