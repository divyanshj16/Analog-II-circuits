*Schmitt Trigger
X1 2 3 4 5 6 ua741
R1 1 3 5k
R2 2 0 10k
R3 2 6 10k
Vcc 4 0 dc 12v
Vee 0 5 dc 12v
Vin 1 0 sin(0 10v 700hz)
.include ua741
.tran 0 10ms 0ms 0.01ms
.probe
.end 
