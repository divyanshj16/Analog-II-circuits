*Square Wave Generator
X1 1 2 3 4 5 ua741
R1 2 5 50
R2 1 0 10k
R3 1 5 1000k
C1 2 0 1mf
Vcc 3 0 dc 12v
Vee 0 4 dc 12v
.include ua741
.tran 0.2us 15ms 5ms 0.001ms
.probe
.end
