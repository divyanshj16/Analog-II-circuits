*Integrator
X1 0 1 3 4 2 ua741
R1 5 1 2k
R2 1 2 24k
C1 1 2 15n
Vcc 3 0 dc 12v
Vee 0 4 dc 12v
Vin 5 0 pulse(0v 1v 0ms 0ms 0ms .1ms .2ms )
.include ua741
.tran .4us 6ms 4ms 0.001ms
.probe
.end
