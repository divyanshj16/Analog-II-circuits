*Non-Inverting Amplifier
x1 1 2 4 5 3 ua741
R1 2 0 1k
Rf 2 3 4k
Vcc 4 0 dc 12v
Vee 0 5 dc 12v
Vin 1 0 sin(0 5mv 1khz)
.include ua741
.tran 0 2ms
.probe
.end
