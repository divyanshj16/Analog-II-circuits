*Peak Detector Circuit
X1 1 2 3 4 5 uA741
D1 0 5 D1N4148
D2 5 6 D1N4148
R1 2 6 10k
R2 1 7 10k
C1 6 0 1n
Vcc 3 0 dc 12v
Vee 0 4 dc 12v
Vin 7 0 sin(0 2v 1khz)
.include ua741
.include D1N4148
.tran 0 2ms
.probe
.end
