*Zero Crossing detector using IC741
X1 1 2 4 5 6 ua741
R1 2 0 1k
R2 1 3 5k
Vin 3 0 sin(0v 5v 50hz 0ms 0hz 0d)
D1 1 2 D1N4148
D2 2 1 D1N4148
Vcc 4 0 dc 12v
Vee 0 5 dc 12v
.include ua741
.include D1N4148
.tran 0 200ms 0ms 200us 
.probe
.end
