*Voltage Follower using Op-Amp
X1 2 1 3 4 1 ua741
Vin 2 0 sin(0 5mv 1khz)
Vcc 3 0 dc 12v
vee 0 4 dc 12v
.include ua741
.tran 0 2ms
.probe
.end


