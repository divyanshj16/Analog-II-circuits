*Precision Rectifier Half Wave
X1 5 2 6 7 3 ua741
D1 2 3 D1N4148
D2 3 4 D1N4148
R1 1 2 10k
R2 2 4 10k
R3 5 0 2k
Vcc 6 0 dc 12v
Vee 0 7 dc 12v
Vin 1 0 sin(0 250mv 1khz)
.include ua741
.include D1N4148
.tran 0 10ms 8ms .001ms
.probe
.end

